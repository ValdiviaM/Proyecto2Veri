
class router_sequence extends uvm_sequence;
	`uvm_object_utils(router_sequence)

endclass:router_sequence
