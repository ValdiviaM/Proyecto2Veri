package pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"


endpackage : pkg    